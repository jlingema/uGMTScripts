

 
 
 

 



window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /virtex7_rx_buf_tb/status
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/CLKA
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/ADDRA
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/DINA
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/WEA
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/CLKB
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/ADDRB
      waveform add -signals /virtex7_rx_buf_tb/virtex7_rx_buf_synth_inst/bmg_port/DOUTB

console submit -using simulator -wait no "run"
